module MIO_BUS( input clk,
			    input rst,
			    input[3:0]BTN,
			    input[15:0]SW,
				
			    input mem_w,
				input mem_r,
			    input[31:0]Cpu_data2bus,				// CPU -> BUS 
			    input[31:0]addr_bus,
			    
				output reg[31:0]Cpu_data4bus,		    // BUS -> CPU
				
				input[31:0]ram_data_out,                // RAM -> BUS data
				
				input[31:0]vram_out,					// VRAM -> BUS data ???RGB???
			    
				input[15:0]led_out,						// led -> BUS
			    
				input[31:0]counter_out,					// counter -> BUS
			    input counter0_out,
			    input counter1_out,
			    input counter2_out,
				
			    input vga_rdn,							// vga -> BUS valid
				
				input ps2_ready,						// ps2 -> BUS valid + pressKey
				input [7:0]key,
				
			    output reg ps2_rdn,						// BUS -> ps2 control/enable
			    
				output reg vram_write,					// BUS -> VRAM control + data + address
			    output reg[11:0]vram_data_in,			// 4R 4G 4B
			    output reg[12:0]cpu_vram_addr,			// cpu write RGB to VRAM
				
				/* VRAM is double port; read/write in different clocks! */
				/* VRAM read address generated by VGAC module  VRAM's data out RGB -> VGAC */
				/* VRAM write address geerate by CPU/BUS; just here! */
				
			    output reg data_ram_we,					// BUS -> RAM control + data + address	 
				output reg[31:0]ram_data_in,			// from CPU write to Memory
				output reg[9:0]ram_addr,				// Memory Address signals
				
			    output reg GPIOffffff00_we,				// BUS -> LED/set control/anable
				
				output reg GPIOfffffe00_we,				// BUS -> segemt control/en
				
			    output reg counter_we,					// BUS -> counter control/en
				
			    output reg[31:0]Peripheral_in 			// BUS -> Peripheral Parallel data except RAM/VRAM
			    );

	wire counter_over;

	//RAM & IO decode signals:	
	always @* begin
		data_ram_we = 0;
		counter_we = 0;
		GPIOffffff00_we = 0;
		GPIOfffffe00_we = 0;
		ram_addr = 10'h0;
		ram_data_in = 32'h0;
		Peripheral_in=32'h0;
		Cpu_data4bus = 32'h0;
		ps2_rdn = 1;
		
		casex(addr_bus[31:8])
			24'h0000xx: begin 				// data_ram (00000000 - 0000ffff(00000ffc), actually lower 4KB RAM)
				data_ram_we = mem_w;
				ram_addr=addr_bus[12:2];   // bit -> word
				ram_data_in=Cpu_data2bus;
				Cpu_data4bus=ram_data_out;			
			end
			24'h000cxx: begin 				// Vram (000c0000 - c000ffff(000012c0), actually lower 4*32KB VRAM)
				vram_write = mem_w ;       // 2^13 = 8 * 1024 = ...
				cpu_vram_addr=addr_bus[12:0];    // just a pixel == just a 12/8 bits == just a row
				vram_data_in=Cpu_data2bus[11:0]; // write vram 8bits / 12bits
				Cpu_data4bus=vga_rdn? {20'h0, vram_out[11:0]} :  32'hx ;			
			end		
			
			24'hffffdx: begin					//PS2 (ffffd000~ ffffdfff)
				ps2_rdn = ~mem_r;
				Peripheral_in = Cpu_data2bus;					    //write NU 
				Cpu_data4bus = {23'h0, ps2_ready, key};				//read from PS2;
			end 

			24'hfffffe: begin  					// 7 Segement LEDs (fffffe00 - fffffeff, 4 7-seg display)
			//24'he00000: begin	
				GPIOfffffe00_we = mem_w;
				Peripheral_in = Cpu_data2bus;
				Cpu_data4bus =counter_out;					//read from Counter
			end
					
			24'hffffff: begin 				  // LED   (ffffff00-ffffffff0,8 LEDs & counter, ffffff04-fffffff4)
			//24'hf00000: begin	
				if(addr_bus[2]) begin		  //ffffff04  for addr of counter
					counter_we = mem_w;
					Peripheral_in = Cpu_data2bus;	    //write Counter Value 
					Cpu_data4bus = counter_out;			//read from Counter;
				end 
				else begin							//ffffff00
					GPIOffffff00_we = mem_w;
					Peripheral_in = Cpu_data2bus;	//write led + 00 counter_set
					//Cpu_data4bus = {counter0_out,counter1_out,counter2_out,17'b0,BTN[3:0],SW[7:0]};
													// read  SW + led_out + counter012_out
					Cpu_data4bus = {counter0_out,counter1_out,counter2_out,led_out[12:0], SW};
				end 
			end
		endcase
	end			// always end

endmodule